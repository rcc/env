library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

--#############################################################################

entity %%% is
    port(
        );  
end entity %%%;

--#############################################################################

architecture RTL of %%% is

    --=========================================================================
    --  Constant declarations
    --=========================================================================



    --=========================================================================
    --  Global Signal declarations
    --=========================================================================



    --=========================================================================
    --  Logic
    --=========================================================================
begin



end architecture RTL;       -- %%%
